module Traffic_Light_Controller (
    input x;
    input clk;
    input clear;
    output reg [1:0] hwy;
    output reg [1:0] cntry;

);
    
endmodule